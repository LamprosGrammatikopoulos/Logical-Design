module f3(x3,b0,b1,b2,b3);
  
	input b0,b1,b2,b3;
	output x3;

       buf gate_buf_1(x3, b0);



endmodule

